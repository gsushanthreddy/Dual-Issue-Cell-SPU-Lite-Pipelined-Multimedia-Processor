package descriptions;
        parameter BYTE = 8;
        parameter HALFWORD = 16;
        parameter WORD = 32;
        parameter QUADWORD = 128;
        parameter ODD = 1;
        parameter EVEN = 0; 

        parameter SMAX = $bitstoshortreal(32'h7fffffff);
        parameter SMIN = $bitstoshortreal(32'h80000000);
        parameter LSLR = 32'h00007FFF;

        typedef enum logic[0:6] {   // logic is defined to handle procedural blocks and continuous assign statements
            ADD_WORD                                                = 7'd1,
            ADD_HALFWORD                                            = 7'd2,
            ADD_HALFWORD_IMMEDIATE                                  = 7'd3,
            ADD_WORD_IMMEDIATE                                      = 7'd4,
            SUBTRACT_FROM_WORD                                      = 7'd5,
            SUBTRACT_FROM_HALFWORD                                  = 7'd6,
            SUBTRACT_FROM_HALFWORD_IMMEDIATE                        = 7'd7,
            SUBTRACT_FROM_WORD_IMMEDIATE                            = 7'd8,
            ADD_EXTENDED                                            = 7'd9,
            SUBTRACT_FROM_EXTENDED                                  = 7'd10,
            CARRY_GENERATE                                          = 7'd11,
            BORROW_GENERATE                                         = 7'd12,
            AND                                                     = 7'd13,
            AND_WITH_COMPLEMENT                                     = 7'd14,
            AND_HALFWORD_IMMEDIATE                                  = 7'd15,
            AND_WORD_IMMEDIATE                                      = 7'd16,
            OR                                                      = 7'd17,
            OR_COMPLEMENT                                           = 7'd18,
            OR_HALFWORD_IMMEDIATE                                   = 7'd19,
            OR_WORD_IMMEDIATE                                       = 7'd20,
            EXCLUSIVE_OR                                            = 7'd21,
            EXCLUSIVE_OR_HALFWORD_IMMEDIATE                         = 7'd22,
            EXCLUSIVE_OR_WORD_IMMEDIATE                             = 7'd23,
            NAND                                                    = 7'd24,
            NOR                                                     = 7'd25,
            COUNT_LEADING_ZEROS                                     = 7'd26,
            FORM_SELECT_MASK_FOR_HALFWORDS                          = 7'd27,
            FORM_SELECT_MASK_FOR_WORDS                              = 7'd28,
            COMPARE_EQUAL_HALFWORD                                  = 7'd29,
            COMPARE_EQUAL_HALFWORD_IMMEDIATE                        = 7'd30,
            COMPARE_EQUAL_WORD                                      = 7'd31,
            COMPARE_EQUAL_WORD_IMMEDIATE                            = 7'd32,
            COMPARE_GREATER_THAN_HALFWORD                           = 7'd33,
            COMPARE_GREATER_THAN_HALFWORD_IMMEDIATE                 = 7'd34,
            COMPARE_GREATER_THAN_WORD                               = 7'd35,
            COMPARE_GREATER_THAN_WORD_IMMEDIATE                     = 7'd36,
            COMPARE_LOGICAL_GREATER_THAN_HALFWORD                   = 7'd37,
            COMPARE_LOGICAL_GREATER_THAN_HALFWORD_IMMEDIATE         = 7'd38,
            COMPARE_LOGICAL_GREATER_THAN_WORD                       = 7'd39,
            COMPARE_LOGICAL_GREATER_THAN_WORD_IMMEDIATE             = 7'd40,
            IMMEDIATE_LOAD_HALFWORD                                 = 7'd41,
            IMMEDIATE_LOAD_HALFWORD_UPPER                           = 7'd42,
            IMMEDIATE_LOAD_WORD                                     = 7'd43,
            IMMEDIATE_LOAD_ADDRESS                                  = 7'd44,
            SHIFT_LEFT_HALFWORD                                     = 7'd45,
            SHIFT_LEFT_HALFWORD_IMMEDIATE                           = 7'd46,
            SHIFT_LEFT_WORD                                         = 7'd47,
            SHIFT_LEFT_WORD_IMMEDIATE                               = 7'd48,
            ROTATE_HALFWORD                                         = 7'd49,
            ROTATE_HALFWORD_IMMEDIATE                               = 7'd50,
            ROTATE_WORD                                             = 7'd51,
            ROTATE_WORD_IMMEDIATE                                   = 7'd52,
            FLOATING_MULTIPLY                                       = 7'd53,
            FLOATING_MULTIPLY_AND_ADD                               = 7'd54,
            FLOATING_NEGATIVE_MULTIPLY_AND_SUBTRACT                 = 7'd55,
            FLOATING_MULTIPLY_AND_SUBTRACT                          = 7'd56,
            MULTIPLY                                                = 7'd57,
            MULTIPLY_UNSIGNED                                       = 7'd58,
            MULTIPLY_IMMEDIATE                                      = 7'd59,
            MULTIPLY_UNSIGNED_IMMEDIATE                             = 7'd60,
            MULTIPLY_AND_ADD                                        = 7'd61,
            MULTIPLY_HIGH                                           = 7'd62,
            ABSOLUTE_DIFFERENCES_OF_BYTES                           = 7'd63,
            AVERAGE_BYTES                                           = 7'd64,
            SUM_BYTES_INTO_HALFWORDS                                = 7'd65,
            COUNT_ONES_IN_BYTES                                     = 7'd66,
            SHIFT_LEFT_QUADWORD_BY_BITS                             = 7'd67,
            SHIFT_LEFT_QUADWORD_BY_BITS_IMMEDIATE                   = 7'd68,
            SHIFT_LEFT_QUADWORD_BY_BYTES                            = 7'd69,
            SHIFT_LEFT_QUADWORD_BY_BYTE_IMMEDIATE                   = 7'd70,
            SHIFT_LEFT_QUADWORD_BY_BYTES_FROM_BIT_SHIFT_COUNT       = 7'd71,
            ROTATE_QUADWORD_BY_BYTES                                = 7'd72,
            ROTATE_QUADWORD_BY_BYTES_IMMEDIATE                      = 7'd73,
            ROTATE_QUADWORD_BY_BYTES_FROM_BIT_SHIFT_COUNT           = 7'd74,
            ROTATE_QUADWORD_BY_BITS                                 = 7'd75,
            ROTATE_QUADWORD_BY_BITS_IMMEDIATE                       = 7'd76,
            GATHER_BITS_FROM_BYTES                                  = 7'd77,
            GATHER_BITS_FROM_HALFWORDS                              = 7'd78,
            GATHER_BITS_FROM_WORDS                                  = 7'd79,
            LOAD_QUADFORM_DFORM                                     = 7'd80,
            LOAD_QUADWORD_AFORM                                     = 7'd81,
            STORE_QUADFORM_DFORM                                    = 7'd82,
            STORE_QUADFORM_AFORM                                    = 7'd83,
            BRANCH_RELATIVE                                         = 7'd84,
            BRANCH_ABSOLUTE                                         = 7'd85,
            BRANCH_RELATIVE_AND_SET_LINK                            = 7'd86,
            BRANCH_ABSOLUTE_AND_SET_LINK                            = 7'd87,
            BRANCH_IF_NOT_ZERO_WORD                                 = 7'd88,
            BRANCH_IF_ZERO_WORD                                     = 7'd89,
            BRANCH_IF_NOT_ZERO_HALFWORD                             = 7'd90,
            BRANCH_IF_ZERO_HALFWORD                                 = 7'd91,
            STOP_AND_SIGNAL                                         = 7'd92,
            NO_OPERATION_EXECUTE                                    = 7'd93,
            NO_OPERATION_LOAD                                       = 7'd94
        } opcode;
endpackage